
`include "opcodes.v"

module control_unit(clk, rst, op,func3, func7 );
    input clk,rst;

    input wire [6:0] op;
    input wire [2:0] func3;
    input wire [6:0] func7;






endmodule